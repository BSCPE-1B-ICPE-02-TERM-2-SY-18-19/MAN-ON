CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 0 1 100 10
342 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
510 176 623 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
2 +V
167 135 282 0 1 3
0 7
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5130 0 0
2
43529 0
0
9 2-In AND~
219 579 241 0 3 22
0 8 4 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
391 0 0
2
43529 0
0
9 2-In AND~
219 437 236 0 3 22
0 6 5 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3124 0 0
2
43529 0
0
7 Ground~
168 987 256 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3421 0 0
2
43529 0
0
9 CC 7-Seg~
183 926 301 0 17 19
10 17 16 15 14 13 12 11 18 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8157 0 0
2
43529 0
0
6 74LS48
188 786 418 0 14 29
0 3 4 5 6 19 20 11 12 13
14 15 16 17 21
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
5572 0 0
2
43529 0
0
6 74112~
219 642 354 0 7 32
0 7 9 10 9 7 22 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8901 0 0
2
43529 0
0
6 74112~
219 498 351 0 7 32
0 7 8 10 8 7 23 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7361 0 0
2
43529 0
0
6 74112~
219 375 351 0 7 32
0 7 6 10 6 7 24 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4747 0 0
2
43529 0
0
6 74112~
219 244 353 0 7 32
0 7 7 10 7 7 25 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
972 0 0
2
43529 0
0
7 Pulser~
4 101 333 0 10 12
0 26 27 10 28 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3472 0 0
2
43529 0
0
36
1 7 3 0 0 16512 0 6 7 0 0 5
754 382
733 382
733 433
666 433
666 318
2 0 4 0 0 12416 0 6 0 0 13 5
754 391
741 391
741 438
531 438
531 315
3 0 5 0 0 12416 0 6 0 0 4 5
754 400
748 400
748 444
403 444
403 315
7 2 5 0 0 0 0 9 3 0 0 3
399 315
413 315
413 245
1 0 6 0 0 4096 0 3 0 0 9 3
413 227
290 227
290 317
4 0 6 0 0 8320 0 6 0 0 9 4
754 409
754 449
272 449
272 317
0 0 7 0 0 4096 0 0 0 23 28 2
283 288
283 373
0 4 6 0 0 0 0 0 9 9 0 3
305 317
305 333
351 333
7 2 6 0 0 0 0 10 9 0 0 4
268 317
337 317
337 315
351 315
0 4 8 0 0 4096 0 0 8 11 0 3
470 315
470 333
474 333
2 0 8 0 0 8192 0 8 0 0 12 3
474 315
464 315
464 236
3 1 8 0 0 4224 0 3 2 0 0 4
458 236
547 236
547 232
555 232
7 2 4 0 0 0 0 8 2 0 0 4
522 315
547 315
547 250
555 250
2 0 9 0 0 4096 0 7 0 0 15 2
618 318
600 318
3 4 9 0 0 4224 0 2 7 0 0 3
600 241
600 336
618 336
4 0 7 0 0 0 0 10 0 0 22 3
220 335
183 335
183 288
3 0 10 0 0 8192 0 10 0 0 20 3
214 326
210 326
210 395
3 0 10 0 0 8192 0 9 0 0 20 3
345 324
341 324
341 395
3 0 10 0 0 0 0 8 0 0 20 3
468 324
464 324
464 395
3 3 10 0 0 12416 0 11 7 0 0 5
125 324
152 324
152 395
612 395
612 327
2 0 7 0 0 0 0 10 0 0 22 3
220 317
210 317
210 288
1 1 7 0 0 8208 0 10 1 0 0 4
244 290
244 288
135 288
135 291
1 1 7 0 0 4096 0 9 10 0 0 3
375 288
244 288
244 290
1 1 7 0 0 0 0 8 9 0 0 2
498 288
375 288
1 1 7 0 0 8192 0 7 8 0 0 3
642 291
642 288
498 288
5 0 7 0 0 0 0 8 0 0 28 3
498 363
498 373
497 373
5 0 7 0 0 0 0 9 0 0 28 2
375 363
375 373
5 5 7 0 0 8320 0 7 10 0 0 4
642 366
642 373
244 373
244 365
7 7 11 0 0 8320 0 5 6 0 0 3
941 337
941 382
818 382
6 8 12 0 0 8320 0 5 6 0 0 3
935 337
935 391
818 391
5 9 13 0 0 8320 0 5 6 0 0 3
929 337
929 400
818 400
4 10 14 0 0 8320 0 5 6 0 0 3
923 337
923 409
818 409
3 11 15 0 0 8320 0 5 6 0 0 3
917 337
917 418
818 418
2 12 16 0 0 8320 0 5 6 0 0 3
911 337
911 427
818 427
13 1 17 0 0 8320 0 6 5 0 0 3
818 436
905 436
905 337
9 1 2 0 0 8320 0 5 4 0 0 4
926 259
926 242
987 242
987 250
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
750 96 883 120
760 104 872 120
14 ______________
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
751 69 884 93
761 77 873 93
14 MARCH 04, 2019
-24 0 0 0 700 0 0 0 0 3 2 1 34
15 Segoe UI Symbol
0 0 0 35
274 136 802 180
284 144 791 176
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
134 94 219 118
144 102 208 118
8 BSCPE-1B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
131 70 296 94
141 78 285 94
18 RAY JOHN J. MAN-ON
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
